--library ieee;
--use ieee.std_logic_1164.all;
--use work.MemoTableTConstants.all;
--
--entity Teste is
----entity Memo_Table_T is 
--	port(
--		--PC address
--		RWAddress: in std_logic_vector(31 downto 0);
--		--Instruction fetched
--		WInstruction: in std_logic_vector(31 downto 0);
--		--Value of the first operand
--		WValue1: in std_logic_vector(31 downto 0);
--		--Value of the second operand
--		WValue2: in std_logic_vector(31 downto 0);
--		--Value of the calculated result
--		WResult: in std_logic_vector(31 downto 0);
--		
--		--Low level activation reset
--		Reset: in std_logic;
--		Clock: in std_logic;
--		
--		--Soltar resultado do ciclo anterior? (Registrador de estado embutido)
--		--Data read from each table way
--		--Data(i)(MemoTableTWidth) = '1' => Hit
--		--Data(i)(MemoTableTWidth) = '0' => Miss
--		
--		Data: out MemoTableTReadData
--	);
----end Memo_Table_T;
--end Teste;
--
----architecture MemoTableTBehaviour of Memo_Table_T is
--architecture MemoTableTBehaviour of Teste is
--
--	
--
--begin
--	
--	
--	
--	process(Clock, Reset)
--	begin
--		
--	end process;
--	
--end MemoTableTBehaviour;