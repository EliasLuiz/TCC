-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: MemoTableTOutput.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any Output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

use work.Constants.all;
use work.DefTypes.all;

ENTITY MemoTableTOutputWay IS
--ENTITY TraceMemory IS
	PORT
	(
		Clock		: IN 	STD_LOGIC  := '1';
		WAddress	: IN 	STD_LOGIC_VECTOR (MemoTableTWayAddressLenght-1 DOWNTO 0);
		WData		: IN 	MemoTableTOutputEntry;
		--WData		: IN 	STD_LOGIC_VECTOR (MemoTableTOutputEntryWidth-1 DOWNTO 0);
		WEnable	: IN 	STD_LOGIC  := '0';
		RAddress	: IN 	STD_LOGIC_VECTOR (MemoTableTWayAddressLenght-1 DOWNTO 0);
		RData		: OUT MemoTableTOutputEntry
		--RData		: OUT STD_LOGIC_VECTOR (MemoTableTOutputEntryWidth-1 DOWNTO 0)
	);
END MemoTableTOutputWay;
--END TraceMemory;


ARCHITECTURE SYN OF MemoTableTOutputWay IS
--ARCHITECTURE SYN OF TraceMemory IS

	SIGNAL RAuxVector : STD_LOGIC_VECTOR (MemoTableTOutputEntryWidth-1 DOWNTO 0);
	SIGNAL WAuxObject : MemoTableTOutputEntry;
	SIGNAL WAuxVector : STD_LOGIC_VECTOR (MemoTableTOutputEntryWidth-1 DOWNTO 0);

	COMPONENT altsyncram
	GENERIC (
		address_reg_b				: STRING;
		clock_enable_input_a		: STRING;
		clock_enable_input_b		: STRING;
		clock_enable_output_a	: STRING;
		clock_enable_output_b	: STRING;
		intended_device_family	: STRING;
		lpm_type						: STRING;
		numwords_a					: NATURAL;
		numwords_b					: NATURAL;
		operation_mode				: STRING;
		outdata_aclr_b				: STRING;
		outdata_reg_b				: STRING;
		power_up_uninitialized	: STRING;
		read_during_write_mode_mixed_ports	: STRING;
		widthad_a			: NATURAL;
		widthad_b			: NATURAL;
		width_a				: NATURAL;
		width_b				: NATURAL;
		width_byteena_a	: NATURAL
	);
	PORT (
		address_a: IN 	STD_LOGIC_VECTOR (MemoTableTWayAddressLenght-1 DOWNTO 0);
		clock0	: IN 	STD_LOGIC;
		data_a	: IN 	STD_LOGIC_VECTOR (MemoTableTOutputEntryWidth-1 DOWNTO 0);
		q_b		: OUT STD_LOGIC_VECTOR (MemoTableTOutputEntryWidth-1 DOWNTO 0);
		wren_a	: IN 	STD_LOGIC;
		address_b: IN 	STD_LOGIC_VECTOR (MemoTableTWayAddressLenght-1 DOWNTO 0)
	);
	END COMPONENT;

BEGIN

	--RData <= RAuxVector;
	RData <= StdLogicToOutput(RAuxVector);
	--WAuxVector <= WData;
	WAuxObject <= WData;
	WAuxVector <= OutputToStdLogic(WAuxObject);

	altsyncram_component : altsyncram
	GENERIC MAP (
		address_reg_b 				=> "CLOCK0",
		clock_enable_input_a 	=> "BYPASS",
		clock_enable_input_b 	=> "BYPASS",
		clock_enable_output_a 	=> "BYPASS",
		clock_enable_output_b 	=> "BYPASS",
		intended_device_family 	=> "Cyclone II",
		lpm_type 					=> "altsyncram",
		numwords_a 					=> MemoTableTWayLenght,
		numwords_b 					=> MemoTableTWayLenght,
		operation_mode 			=> "DUAL_PORT",
		outdata_aclr_b 			=> "NONE",
		outdata_reg_b 				=> "CLOCK0",
		power_up_uninitialized 	=> "FALSE",
		read_during_write_mode_mixed_ports => "DONT_CARE",
		widthad_a 			=> MemoTableTWayAddressLenght,
		widthad_b 			=> MemoTableTWayAddressLenght,
		width_a 				=> MemoTableTOutputEntryWidth,
		width_b 				=> MemoTableTOutputEntryWidth,
		width_byteena_a 	=> 1
	)
	PORT MAP (
		address_a => WAddress,
		clock0 	 => Clock,
		data_a 	 => WAuxVector,
		wren_a 	 => WEnable,
		address_b => RAddress,
		q_b 		 => RAuxVector
	);


END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: ADDRESSSTALL_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_B NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_Output_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_Output_B NUMERIC "0"
-- Retrieval info: PRIVATE: CLRdata NUMERIC "0"
-- Retrieval info: PRIVATE: CLRq NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrdaddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrren NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwraddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwren NUMERIC "0"
-- Retrieval info: PRIVATE: Clock NUMERIC "0"
-- Retrieval info: PRIVATE: Clock_A NUMERIC "0"
-- Retrieval info: PRIVATE: Clock_B NUMERIC "0"
-- Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_REG_B NUMERIC "0"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_B"
-- Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MEMSIZE NUMERIC "4096"
-- Retrieval info: PRIVATE: MEM_IN_BITS NUMERIC "1"
-- Retrieval info: PRIVATE: MIFfilename STRING ""
-- Retrieval info: PRIVATE: OPERATION_MODE NUMERIC "2"
-- Retrieval info: PRIVATE: OUTDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: OUTDATA_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_MIXED_PORTS NUMERIC "2"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_B NUMERIC "3"
-- Retrieval info: PRIVATE: REGdata NUMERIC "1"
-- Retrieval info: PRIVATE: REGq NUMERIC "1"
-- Retrieval info: PRIVATE: REGrdaddress NUMERIC "1"
-- Retrieval info: PRIVATE: REGrren NUMERIC "1"
-- Retrieval info: PRIVATE: REGwraddress NUMERIC "1"
-- Retrieval info: PRIVATE: REGwren NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "1"
-- Retrieval info: PRIVATE: USE_DIFF_CLKEN NUMERIC "0"
-- Retrieval info: PRIVATE: UseDPRAM NUMERIC "1"
-- Retrieval info: PRIVATE: VarWidth NUMERIC "0"
-- Retrieval info: PRIVATE: WIDTH_READ_A NUMERIC "64"
-- Retrieval info: PRIVATE: WIDTH_READ_B NUMERIC "64"
-- Retrieval info: PRIVATE: WIDTH_WRITE_A NUMERIC "64"
-- Retrieval info: PRIVATE: WIDTH_WRITE_B NUMERIC "64"
-- Retrieval info: PRIVATE: WRADDR_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: WRADDR_REG_B NUMERIC "0"
-- Retrieval info: PRIVATE: WRCTRL_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: enable NUMERIC "0"
-- Retrieval info: PRIVATE: rden NUMERIC "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ADDRESS_REG_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_B STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_Output_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_Output_B STRING "BYPASS"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "64"
-- Retrieval info: CONSTANT: NUMWORDS_B NUMERIC "64"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "DUAL_PORT"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_REG_B STRING "CLOCK0"
-- Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_MIXED_PORTS STRING "DONT_CARE"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "6"
-- Retrieval info: CONSTANT: WIDTHAD_B NUMERIC "6"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "64"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "64"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
-- Retrieval info: USED_PORT: data 0 0 64 0 INPUT NODEFVAL "data[MemoTableTOutputEntryWidth-1..0]"
-- Retrieval info: USED_PORT: q 0 0 64 0 Output NODEFVAL "q[MemoTableTOutputEntryWidth-1..0]"
-- Retrieval info: USED_PORT: rdaddress 0 0 6 0 INPUT NODEFVAL "rdaddress[MemoTableTWayAddressLenght-1..0]"
-- Retrieval info: USED_PORT: wraddress 0 0 6 0 INPUT NODEFVAL "wraddress[MemoTableTWayAddressLenght-1..0]"
-- Retrieval info: USED_PORT: wren 0 0 0 0 INPUT GND "wren"
-- Retrieval info: CONNECT: @address_a 0 0 6 0 wraddress 0 0 6 0
-- Retrieval info: CONNECT: @address_b 0 0 6 0 rdaddress 0 0 6 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data_a 0 0 64 0 data 0 0 64 0
-- Retrieval info: CONNECT: @wren_a 0 0 0 0 wren 0 0 0 0
-- Retrieval info: CONNECT: q 0 0 64 0 @q_b 0 0 64 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL MemoTableTOutput.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MemoTableTOutput.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MemoTableTOutput.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MemoTableTOutput.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MemoTableTOutput_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL MemoTableTOutput_syn.v TRUE
-- Retrieval info: LIB_FILE: altera_mf
